package csr_ids_pkg;
  // csr id enum
  import cosim_constants_pkg::REG_KEY_ID_W;
  
  // riscv-isa-sim/riscv/encoding.h dosyasindan
  typedef enum bit unsigned [REG_KEY_ID_W-1:0] {
    CSR_FFLAGS         =  'h1,
    CSR_FRM            =  'h2,
    CSR_FCSR           =  'h3,
    CSR_VSTART         =  'h8,
    CSR_VXSAT          =  'h9,
    CSR_VXRM           =  'ha,
    CSR_VCSR           =  'hf,
    CSR_SEED           =  'h15,
    CSR_JVT            =  'h17,
    CSR_CYCLE          =  'hc00,
    CSR_TIME           =  'hc01,
    CSR_INSTRET        =  'hc02,
    CSR_HPMCOUNTER3    =  'hc03,
    CSR_HPMCOUNTER4    =  'hc04,
    CSR_HPMCOUNTER5    =  'hc05,
    CSR_HPMCOUNTER6    =  'hc06,
    CSR_HPMCOUNTER7    =  'hc07,
    CSR_HPMCOUNTER8    =  'hc08,
    CSR_HPMCOUNTER9    =  'hc09,
    CSR_HPMCOUNTER10   =  'hc0a,
    CSR_HPMCOUNTER11   =  'hc0b,
    CSR_HPMCOUNTER12   =  'hc0c,
    CSR_HPMCOUNTER13   =  'hc0d,
    CSR_HPMCOUNTER14   =  'hc0e,
    CSR_HPMCOUNTER15   =  'hc0f,
    CSR_HPMCOUNTER16   =  'hc10,
    CSR_HPMCOUNTER17   =  'hc11,
    CSR_HPMCOUNTER18   =  'hc12,
    CSR_HPMCOUNTER19   =  'hc13,
    CSR_HPMCOUNTER20   =  'hc14,
    CSR_HPMCOUNTER21   =  'hc15,
    CSR_HPMCOUNTER22   =  'hc16,
    CSR_HPMCOUNTER23   =  'hc17,
    CSR_HPMCOUNTER24   =  'hc18,
    CSR_HPMCOUNTER25   =  'hc19,
    CSR_HPMCOUNTER26   =  'hc1a,
    CSR_HPMCOUNTER27   =  'hc1b,
    CSR_HPMCOUNTER28   =  'hc1c,
    CSR_HPMCOUNTER29   =  'hc1d,
    CSR_HPMCOUNTER30   =  'hc1e,
    CSR_HPMCOUNTER31   =  'hc1f,
    CSR_VL             =  'hc20,
    CSR_VTYPE          =  'hc21,
    CSR_VLENB          =  'hc22,
    CSR_SSTATUS        =  'h100,
    CSR_SEDELEG        =  'h102,
    CSR_SIDELEG        =  'h103,
    CSR_SIE            =  'h104,
    CSR_STVEC          =  'h105,
    CSR_SCOUNTEREN     =  'h106,
    CSR_SENVCFG        =  'h10a,
    CSR_SSTATEEN0      =  'h10c,
    CSR_SSTATEEN1      =  'h10d,
    CSR_SSTATEEN2      =  'h10e,
    CSR_SSTATEEN3      =  'h10f,
    CSR_SCOUNTINHIBIT  =  'h120,
    CSR_SSCRATCH       =  'h140,
    CSR_SEPC           =  'h141,
    CSR_SCAUSE         =  'h142,
    CSR_STVAL          =  'h143,
    CSR_SIP            =  'h144,
    CSR_STIMECMP       =  'h14d,
    CSR_SISELECT       =  'h150,
    CSR_SIREG          =  'h151,
    CSR_SIREG2         =  'h152,
    CSR_SIREG3         =  'h153,
    CSR_SIREG4         =  'h155,
    CSR_SIREG5         =  'h156,
    CSR_SIREG6         =  'h157,
    CSR_STOPEI         =  'h15c,
    CSR_SATP           =  'h180,
    CSR_SCONTEXT       =  'h5a8,
    CSR_VSSTATUS       =  'h200,
    CSR_VSIE           =  'h204,
    CSR_VSTVEC         =  'h205,
    CSR_VSSCRATCH      =  'h240,
    CSR_VSEPC          =  'h241,
    CSR_VSCAUSE        =  'h242,
    CSR_VSTVAL         =  'h243,
    CSR_VSIP           =  'h244,
    CSR_VSTIMECMP      =  'h24d,
    CSR_VSISELECT      =  'h250,
    CSR_VSIREG         =  'h251,
    CSR_VSIREG2        =  'h252,
    CSR_VSIREG3        =  'h253,
    CSR_VSIREG4        =  'h255,
    CSR_VSIREG5        =  'h256,
    CSR_VSIREG6        =  'h257,
    CSR_VSTOPEI        =  'h25c,
    CSR_VSATP          =  'h280,
    CSR_HSTATUS        =  'h600,
    CSR_HEDELEG        =  'h602,
    CSR_HIDELEG        =  'h603,
    CSR_HIE            =  'h604,
    CSR_HTIMEDELTA     =  'h605,
    CSR_HCOUNTEREN     =  'h606,
    CSR_HGEIE          =  'h607,
    CSR_HVIEN          =  'h608,
    CSR_HVICTL         =  'h609,
    CSR_HENVCFG        =  'h60a,
    CSR_HSTATEEN0      =  'h60c,
    CSR_HSTATEEN1      =  'h60d,
    CSR_HSTATEEN2      =  'h60e,
    CSR_HSTATEEN3      =  'h60f,
    CSR_HTVAL          =  'h643,
    CSR_HIP            =  'h644,
    CSR_HVIP           =  'h645,
    CSR_HVIPRIO1       =  'h646,
    CSR_HVIPRIO2       =  'h647,
    CSR_HTINST         =  'h64a,
    CSR_HGATP          =  'h680,
    CSR_HCONTEXT       =  'h6a8,
    CSR_HGEIP          =  'he12,
    CSR_VSTOPI         =  'heb0,
    CSR_SCOUNTOVF      =  'hda0,
    CSR_STOPI          =  'hdb0,
    CSR_UTVT           =  'h7,
    CSR_UNXTI          =  'h45,
    CSR_UINTSTATUS     =  'h46,
    CSR_USCRATCHCSW    =  'h48,
    CSR_USCRATCHCSWL   =  'h49,
    CSR_STVT           =  'h107,
    CSR_SNXTI          =  'h145,
    CSR_SINTSTATUS     =  'h146,
    CSR_SSCRATCHCSW    =  'h148,
    CSR_SSCRATCHCSWL   =  'h149,
    CSR_MTVT           =  'h307,
    CSR_MNXTI          =  'h345,
    CSR_MINTSTATUS     =  'h346,
    CSR_MSCRATCHCSW    =  'h348,
    CSR_MSCRATCHCSWL   =  'h349,
    CSR_MSTATUS        =  'h300,
    CSR_MISA           =  'h301,
    CSR_MEDELEG        =  'h302,
    CSR_MIDELEG        =  'h303,
    CSR_MIE            =  'h304,
    CSR_MTVEC          =  'h305,
    CSR_MCOUNTEREN     =  'h306,
    CSR_MVIEN          =  'h308,
    CSR_MVIP           =  'h309,
    CSR_MENVCFG        =  'h30a,
    CSR_MSTATEEN0      =  'h30c,
    CSR_MSTATEEN1      =  'h30d,
    CSR_MSTATEEN2      =  'h30e,
    CSR_MSTATEEN3      =  'h30f,
    CSR_MCOUNTINHIBIT  =  'h320,
    CSR_MSCRATCH       =  'h340,
    CSR_MEPC           =  'h341,
    CSR_MCAUSE         =  'h342,
    CSR_MTVAL          =  'h343,
    CSR_MIP            =  'h344,
    CSR_MTINST         =  'h34a,
    CSR_MTVAL2         =  'h34b,
    CSR_MISELECT       =  'h350,
    CSR_MIREG          =  'h351,
    CSR_MIREG2         =  'h352,
    CSR_MIREG3         =  'h353,
    CSR_MIREG4         =  'h355,
    CSR_MIREG5         =  'h356,
    CSR_MIREG6         =  'h357,
    CSR_MTOPEI         =  'h35c,
    CSR_PMPCFG0        =  'h3a0,
    CSR_PMPCFG1        =  'h3a1,
    CSR_PMPCFG2        =  'h3a2,
    CSR_PMPCFG3        =  'h3a3,
    CSR_PMPCFG4        =  'h3a4,
    CSR_PMPCFG5        =  'h3a5,
    CSR_PMPCFG6        =  'h3a6,
    CSR_PMPCFG7        =  'h3a7,
    CSR_PMPCFG8        =  'h3a8,
    CSR_PMPCFG9        =  'h3a9,
    CSR_PMPCFG10       =  'h3aa,
    CSR_PMPCFG11       =  'h3ab,
    CSR_PMPCFG12       =  'h3ac,
    CSR_PMPCFG13       =  'h3ad,
    CSR_PMPCFG14       =  'h3ae,
    CSR_PMPCFG15       =  'h3af,
    CSR_PMPADDR0       =  'h3b0,
    CSR_PMPADDR1       =  'h3b1,
    CSR_PMPADDR2       =  'h3b2,
    CSR_PMPADDR3       =  'h3b3,
    CSR_PMPADDR4       =  'h3b4,
    CSR_PMPADDR5       =  'h3b5,
    CSR_PMPADDR6       =  'h3b6,
    CSR_PMPADDR7       =  'h3b7,
    CSR_PMPADDR8       =  'h3b8,
    CSR_PMPADDR9       =  'h3b9,
    CSR_PMPADDR10      =  'h3ba,
    CSR_PMPADDR11      =  'h3bb,
    CSR_PMPADDR12      =  'h3bc,
    CSR_PMPADDR13      =  'h3bd,
    CSR_PMPADDR14      =  'h3be,
    CSR_PMPADDR15      =  'h3bf,
    CSR_PMPADDR16      =  'h3c0,
    CSR_PMPADDR17      =  'h3c1,
    CSR_PMPADDR18      =  'h3c2,
    CSR_PMPADDR19      =  'h3c3,
    CSR_PMPADDR20      =  'h3c4,
    CSR_PMPADDR21      =  'h3c5,
    CSR_PMPADDR22      =  'h3c6,
    CSR_PMPADDR23      =  'h3c7,
    CSR_PMPADDR24      =  'h3c8,
    CSR_PMPADDR25      =  'h3c9,
    CSR_PMPADDR26      =  'h3ca,
    CSR_PMPADDR27      =  'h3cb,
    CSR_PMPADDR28      =  'h3cc,
    CSR_PMPADDR29      =  'h3cd,
    CSR_PMPADDR30      =  'h3ce,
    CSR_PMPADDR31      =  'h3cf,
    CSR_PMPADDR32      =  'h3d0,
    CSR_PMPADDR33      =  'h3d1,
    CSR_PMPADDR34      =  'h3d2,
    CSR_PMPADDR35      =  'h3d3,
    CSR_PMPADDR36      =  'h3d4,
    CSR_PMPADDR37      =  'h3d5,
    CSR_PMPADDR38      =  'h3d6,
    CSR_PMPADDR39      =  'h3d7,
    CSR_PMPADDR40      =  'h3d8,
    CSR_PMPADDR41      =  'h3d9,
    CSR_PMPADDR42      =  'h3da,
    CSR_PMPADDR43      =  'h3db,
    CSR_PMPADDR44      =  'h3dc,
    CSR_PMPADDR45      =  'h3dd,
    CSR_PMPADDR46      =  'h3de,
    CSR_PMPADDR47      =  'h3df,
    CSR_PMPADDR48      =  'h3e0,
    CSR_PMPADDR49      =  'h3e1,
    CSR_PMPADDR50      =  'h3e2,
    CSR_PMPADDR51      =  'h3e3,
    CSR_PMPADDR52      =  'h3e4,
    CSR_PMPADDR53      =  'h3e5,
    CSR_PMPADDR54      =  'h3e6,
    CSR_PMPADDR55      =  'h3e7,
    CSR_PMPADDR56      =  'h3e8,
    CSR_PMPADDR57      =  'h3e9,
    CSR_PMPADDR58      =  'h3ea,
    CSR_PMPADDR59      =  'h3eb,
    CSR_PMPADDR60      =  'h3ec,
    CSR_PMPADDR61      =  'h3ed,
    CSR_PMPADDR62      =  'h3ee,
    CSR_PMPADDR63      =  'h3ef,
    CSR_MSECCFG        =  'h747,
    CSR_TSELECT        =  'h7a0,
    CSR_TDATA1         =  'h7a1,
    CSR_TDATA2         =  'h7a2,
    CSR_TDATA3         =  'h7a3,
    CSR_TINFO          =  'h7a4,
    CSR_TCONTROL       =  'h7a5,
    CSR_MCONTEXT       =  'h7a8,
    CSR_MSCONTEXT      =  'h7aa,
    CSR_DCSR           =  'h7b0,
    CSR_DPC            =  'h7b1,
    CSR_DSCRATCH0      =  'h7b2,
    CSR_DSCRATCH1      =  'h7b3,
    CSR_MCYCLE         =  'hb00,
    CSR_MINSTRET       =  'hb02,
    CSR_MHPMCOUNTER3   =  'hb03,
    CSR_MHPMCOUNTER4   =  'hb04,
    CSR_MHPMCOUNTER5   =  'hb05,
    CSR_MHPMCOUNTER6   =  'hb06,
    CSR_MHPMCOUNTER7   =  'hb07,
    CSR_MHPMCOUNTER8   =  'hb08,
    CSR_MHPMCOUNTER9   =  'hb09,
    CSR_MHPMCOUNTER10  =  'hb0a,
    CSR_MHPMCOUNTER11  =  'hb0b,
    CSR_MHPMCOUNTER12  =  'hb0c,
    CSR_MHPMCOUNTER13  =  'hb0d,
    CSR_MHPMCOUNTER14  =  'hb0e,
    CSR_MHPMCOUNTER15  =  'hb0f,
    CSR_MHPMCOUNTER16  =  'hb10,
    CSR_MHPMCOUNTER17  =  'hb11,
    CSR_MHPMCOUNTER18  =  'hb12,
    CSR_MHPMCOUNTER19  =  'hb13,
    CSR_MHPMCOUNTER20  =  'hb14,
    CSR_MHPMCOUNTER21  =  'hb15,
    CSR_MHPMCOUNTER22  =  'hb16,
    CSR_MHPMCOUNTER23  =  'hb17,
    CSR_MHPMCOUNTER24  =  'hb18,
    CSR_MHPMCOUNTER25  =  'hb19,
    CSR_MHPMCOUNTER26  =  'hb1a,
    CSR_MHPMCOUNTER27  =  'hb1b,
    CSR_MHPMCOUNTER28  =  'hb1c,
    CSR_MHPMCOUNTER29  =  'hb1d,
    CSR_MHPMCOUNTER30  =  'hb1e,
    CSR_MHPMCOUNTER31  =  'hb1f,
    CSR_MCYCLECFG      =  'h321,
    CSR_MINSTRETCFG    =  'h322,
    CSR_MHPMEVENT3     =  'h323,
    CSR_MHPMEVENT4     =  'h324,
    CSR_MHPMEVENT5     =  'h325,
    CSR_MHPMEVENT6     =  'h326,
    CSR_MHPMEVENT7     =  'h327,
    CSR_MHPMEVENT8     =  'h328,
    CSR_MHPMEVENT9     =  'h329,
    CSR_MHPMEVENT10    =  'h32a,
    CSR_MHPMEVENT11    =  'h32b,
    CSR_MHPMEVENT12    =  'h32c,
    CSR_MHPMEVENT13    =  'h32d,
    CSR_MHPMEVENT14    =  'h32e,
    CSR_MHPMEVENT15    =  'h32f,
    CSR_MHPMEVENT16    =  'h330,
    CSR_MHPMEVENT17    =  'h331,
    CSR_MHPMEVENT18    =  'h332,
    CSR_MHPMEVENT19    =  'h333,
    CSR_MHPMEVENT20    =  'h334,
    CSR_MHPMEVENT21    =  'h335,
    CSR_MHPMEVENT22    =  'h336,
    CSR_MHPMEVENT23    =  'h337,
    CSR_MHPMEVENT24    =  'h338,
    CSR_MHPMEVENT25    =  'h339,
    CSR_MHPMEVENT26    =  'h33a,
    CSR_MHPMEVENT27    =  'h33b,
    CSR_MHPMEVENT28    =  'h33c,
    CSR_MHPMEVENT29    =  'h33d,
    CSR_MHPMEVENT30    =  'h33e,
    CSR_MHPMEVENT31    =  'h33f,
    CSR_MVENDORID      =  'hf11,
    CSR_MARCHID        =  'hf12,
    CSR_MIMPID         =  'hf13,
    CSR_MHARTID        =  'hf14,
    CSR_MCONFIGPTR     =  'hf15,
    CSR_MTOPI          =  'hfb0,
    CSR_SIEH           =  'h114,
    CSR_SIPH           =  'h154,
    CSR_STIMECMPH      =  'h15d,
    CSR_VSIEH          =  'h214,
    CSR_VSIPH          =  'h254,
    CSR_VSTIMECMPH     =  'h25d,
    CSR_HTIMEDELTAH    =  'h615,
    CSR_HIDELEGH       =  'h613,
    CSR_HVIENH         =  'h618,
    CSR_HENVCFGH       =  'h61a,
    CSR_HVIPH          =  'h655,
    CSR_HVIPRIO1H      =  'h656,
    CSR_HVIPRIO2H      =  'h657,
    CSR_HSTATEEN0H     =  'h61c,
    CSR_HSTATEEN1H     =  'h61d,
    CSR_HSTATEEN2H     =  'h61e,
    CSR_HSTATEEN3H     =  'h61f,
    CSR_CYCLEH         =  'hc80,
    CSR_TIMEH          =  'hc81,
    CSR_INSTRETH       =  'hc82,
    CSR_HPMCOUNTER3H   =  'hc83,
    CSR_HPMCOUNTER4H   =  'hc84,
    CSR_HPMCOUNTER5H   =  'hc85,
    CSR_HPMCOUNTER6H   =  'hc86,
    CSR_HPMCOUNTER7H   =  'hc87,
    CSR_HPMCOUNTER8H   =  'hc88,
    CSR_HPMCOUNTER9H   =  'hc89,
    CSR_HPMCOUNTER10H  =  'hc8a,
    CSR_HPMCOUNTER11H  =  'hc8b,
    CSR_HPMCOUNTER12H  =  'hc8c,
    CSR_HPMCOUNTER13H  =  'hc8d,
    CSR_HPMCOUNTER14H  =  'hc8e,
    CSR_HPMCOUNTER15H  =  'hc8f,
    CSR_HPMCOUNTER16H  =  'hc90,
    CSR_HPMCOUNTER17H  =  'hc91,
    CSR_HPMCOUNTER18H  =  'hc92,
    CSR_HPMCOUNTER19H  =  'hc93,
    CSR_HPMCOUNTER20H  =  'hc94,
    CSR_HPMCOUNTER21H  =  'hc95,
    CSR_HPMCOUNTER22H  =  'hc96,
    CSR_HPMCOUNTER23H  =  'hc97,
    CSR_HPMCOUNTER24H  =  'hc98,
    CSR_HPMCOUNTER25H  =  'hc99,
    CSR_HPMCOUNTER26H  =  'hc9a,
    CSR_HPMCOUNTER27H  =  'hc9b,
    CSR_HPMCOUNTER28H  =  'hc9c,
    CSR_HPMCOUNTER29H  =  'hc9d,
    CSR_HPMCOUNTER30H  =  'hc9e,
    CSR_HPMCOUNTER31H  =  'hc9f,
    CSR_MSTATUSH       =  'h310,
    CSR_MIDELEGH       =  'h313,
    CSR_MIEH           =  'h314,
    CSR_MVIENH         =  'h318,
    CSR_MVIPH          =  'h319,
    CSR_MENVCFGH       =  'h31a,
    CSR_MSTATEEN0H     =  'h31c,
    CSR_MSTATEEN1H     =  'h31d,
    CSR_MSTATEEN2H     =  'h31e,
    CSR_MSTATEEN3H     =  'h31f,
    CSR_MIPH           =  'h354,
    CSR_MCYCLECFGH     =  'h721,
    CSR_MINSTRETCFGH   =  'h722,
    CSR_MHPMEVENT3H    =  'h723,
    CSR_MHPMEVENT4H    =  'h724,
    CSR_MHPMEVENT5H    =  'h725,
    CSR_MHPMEVENT6H    =  'h726,
    CSR_MHPMEVENT7H    =  'h727,
    CSR_MHPMEVENT8H    =  'h728,
    CSR_MHPMEVENT9H    =  'h729,
    CSR_MHPMEVENT10H   =  'h72a,
    CSR_MHPMEVENT11H   =  'h72b,
    CSR_MHPMEVENT12H   =  'h72c,
    CSR_MHPMEVENT13H   =  'h72d,
    CSR_MHPMEVENT14H   =  'h72e,
    CSR_MHPMEVENT15H   =  'h72f,
    CSR_MHPMEVENT16H   =  'h730,
    CSR_MHPMEVENT17H   =  'h731,
    CSR_MHPMEVENT18H   =  'h732,
    CSR_MHPMEVENT19H   =  'h733,
    CSR_MHPMEVENT20H   =  'h734,
    CSR_MHPMEVENT21H   =  'h735,
    CSR_MHPMEVENT22H   =  'h736,
    CSR_MHPMEVENT23H   =  'h737,
    CSR_MHPMEVENT24H   =  'h738,
    CSR_MHPMEVENT25H   =  'h739,
    CSR_MHPMEVENT26H   =  'h73a,
    CSR_MHPMEVENT27H   =  'h73b,
    CSR_MHPMEVENT28H   =  'h73c,
    CSR_MHPMEVENT29H   =  'h73d,
    CSR_MHPMEVENT30H   =  'h73e,
    CSR_MHPMEVENT31H   =  'h73f,
    CSR_MNSCRATCH      =  'h740,
    CSR_MNEPC          =  'h741,
    CSR_MNCAUSE        =  'h742,
    CSR_MNSTATUS       =  'h744,
    CSR_MSECCFGH       =  'h757,
    CSR_MCYCLEH        =  'hb80,
    CSR_MINSTRETH      =  'hb82,
    CSR_MHPMCOUNTER3H  =  'hb83,
    CSR_MHPMCOUNTER4H  =  'hb84,
    CSR_MHPMCOUNTER5H  =  'hb85,
    CSR_MHPMCOUNTER6H  =  'hb86,
    CSR_MHPMCOUNTER7H  =  'hb87,
    CSR_MHPMCOUNTER8H  =  'hb88,
    CSR_MHPMCOUNTER9H  =  'hb89,
    CSR_MHPMCOUNTER10H =  'hb8a,
    CSR_MHPMCOUNTER11H =  'hb8b,
    CSR_MHPMCOUNTER12H =  'hb8c,
    CSR_MHPMCOUNTER13H =  'hb8d,
    CSR_MHPMCOUNTER14H =  'hb8e,
    CSR_MHPMCOUNTER15H =  'hb8f,
    CSR_MHPMCOUNTER16H =  'hb90,
    CSR_MHPMCOUNTER17H =  'hb91,
    CSR_MHPMCOUNTER18H =  'hb92,
    CSR_MHPMCOUNTER19H =  'hb93,
    CSR_MHPMCOUNTER20H =  'hb94,
    CSR_MHPMCOUNTER21H =  'hb95,
    CSR_MHPMCOUNTER22H =  'hb96,
    CSR_MHPMCOUNTER23H =  'hb97,
    CSR_MHPMCOUNTER24H =  'hb98,
    CSR_MHPMCOUNTER25H =  'hb99,
    CSR_MHPMCOUNTER26H =  'hb9a,
    CSR_MHPMCOUNTER27H =  'hb9b,
    CSR_MHPMCOUNTER28H =  'hb9c,
    CSR_MHPMCOUNTER29H =  'hb9d,
    CSR_MHPMCOUNTER30H =  'hb9e,
    CSR_MHPMCOUNTER31H =  'hb9f
  } csr_id_e;
endpackage