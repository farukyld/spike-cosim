package csr_ids_pkg;
  // csr id enum
  import cosim_constants_pkg::REG_KEY_ID_W;
  typedef enum bit [REG_KEY_ID_W-1:0] {
    // riscv/encoding.h
    CSR_FFLAGS         =  REG_KEY_ID_W'('h1),
    CSR_FRM            =  REG_KEY_ID_W'('h2),
    CSR_FCSR           =  REG_KEY_ID_W'('h3),
    CSR_VSTART         =  REG_KEY_ID_W'('h8),
    CSR_VXSAT          =  REG_KEY_ID_W'('h9),
    CSR_VXRM           =  REG_KEY_ID_W'('ha),
    CSR_VCSR           =  REG_KEY_ID_W'('hf),
    CSR_SEED           =  REG_KEY_ID_W'('h15),
    CSR_JVT            =  REG_KEY_ID_W'('h17),
    CSR_CYCLE          =  REG_KEY_ID_W'('hc00),
    CSR_TIME           =  REG_KEY_ID_W'('hc01),
    CSR_INSTRET        =  REG_KEY_ID_W'('hc02),
    CSR_HPMCOUNTER3    =  REG_KEY_ID_W'('hc03),
    CSR_HPMCOUNTER4    =  REG_KEY_ID_W'('hc04),
    CSR_HPMCOUNTER5    =  REG_KEY_ID_W'('hc05),
    CSR_HPMCOUNTER6    =  REG_KEY_ID_W'('hc06),
    CSR_HPMCOUNTER7    =  REG_KEY_ID_W'('hc07),
    CSR_HPMCOUNTER8    =  REG_KEY_ID_W'('hc08),
    CSR_HPMCOUNTER9    =  REG_KEY_ID_W'('hc09),
    CSR_HPMCOUNTER10   =  REG_KEY_ID_W'('hc0a),
    CSR_HPMCOUNTER11   =  REG_KEY_ID_W'('hc0b),
    CSR_HPMCOUNTER12   =  REG_KEY_ID_W'('hc0c),
    CSR_HPMCOUNTER13   =  REG_KEY_ID_W'('hc0d),
    CSR_HPMCOUNTER14   =  REG_KEY_ID_W'('hc0e),
    CSR_HPMCOUNTER15   =  REG_KEY_ID_W'('hc0f),
    CSR_HPMCOUNTER16   =  REG_KEY_ID_W'('hc10),
    CSR_HPMCOUNTER17   =  REG_KEY_ID_W'('hc11),
    CSR_HPMCOUNTER18   =  REG_KEY_ID_W'('hc12),
    CSR_HPMCOUNTER19   =  REG_KEY_ID_W'('hc13),
    CSR_HPMCOUNTER20   =  REG_KEY_ID_W'('hc14),
    CSR_HPMCOUNTER21   =  REG_KEY_ID_W'('hc15),
    CSR_HPMCOUNTER22   =  REG_KEY_ID_W'('hc16),
    CSR_HPMCOUNTER23   =  REG_KEY_ID_W'('hc17),
    CSR_HPMCOUNTER24   =  REG_KEY_ID_W'('hc18),
    CSR_HPMCOUNTER25   =  REG_KEY_ID_W'('hc19),
    CSR_HPMCOUNTER26   =  REG_KEY_ID_W'('hc1a),
    CSR_HPMCOUNTER27   =  REG_KEY_ID_W'('hc1b),
    CSR_HPMCOUNTER28   =  REG_KEY_ID_W'('hc1c),
    CSR_HPMCOUNTER29   =  REG_KEY_ID_W'('hc1d),
    CSR_HPMCOUNTER30   =  REG_KEY_ID_W'('hc1e),
    CSR_HPMCOUNTER31   =  REG_KEY_ID_W'('hc1f),
    CSR_VL             =  REG_KEY_ID_W'('hc20),
    CSR_VTYPE          =  REG_KEY_ID_W'('hc21),
    CSR_VLENB          =  REG_KEY_ID_W'('hc22),
    CSR_SSTATUS        =  REG_KEY_ID_W'('h100),
    CSR_SEDELEG        =  REG_KEY_ID_W'('h102),
    CSR_SIDELEG        =  REG_KEY_ID_W'('h103),
    CSR_SIE            =  REG_KEY_ID_W'('h104),
    CSR_STVEC          =  REG_KEY_ID_W'('h105),
    CSR_SCOUNTEREN     =  REG_KEY_ID_W'('h106),
    CSR_SENVCFG        =  REG_KEY_ID_W'('h10a),
    CSR_SSTATEEN0      =  REG_KEY_ID_W'('h10c),
    CSR_SSTATEEN1      =  REG_KEY_ID_W'('h10d),
    CSR_SSTATEEN2      =  REG_KEY_ID_W'('h10e),
    CSR_SSTATEEN3      =  REG_KEY_ID_W'('h10f),
    CSR_SCOUNTINHIBIT  =  REG_KEY_ID_W'('h120),
    CSR_SSCRATCH       =  REG_KEY_ID_W'('h140),
    CSR_SEPC           =  REG_KEY_ID_W'('h141),
    CSR_SCAUSE         =  REG_KEY_ID_W'('h142),
    CSR_STVAL          =  REG_KEY_ID_W'('h143),
    CSR_SIP            =  REG_KEY_ID_W'('h144),
    CSR_STIMECMP       =  REG_KEY_ID_W'('h14d),
    CSR_SISELECT       =  REG_KEY_ID_W'('h150),
    CSR_SIREG          =  REG_KEY_ID_W'('h151),
    CSR_SIREG2         =  REG_KEY_ID_W'('h152),
    CSR_SIREG3         =  REG_KEY_ID_W'('h153),
    CSR_SIREG4         =  REG_KEY_ID_W'('h155),
    CSR_SIREG5         =  REG_KEY_ID_W'('h156),
    CSR_SIREG6         =  REG_KEY_ID_W'('h157),
    CSR_STOPEI         =  REG_KEY_ID_W'('h15c),
    CSR_SATP           =  REG_KEY_ID_W'('h180),
    CSR_SCONTEXT       =  REG_KEY_ID_W'('h5a8),
    CSR_VSSTATUS       =  REG_KEY_ID_W'('h200),
    CSR_VSIE           =  REG_KEY_ID_W'('h204),
    CSR_VSTVEC         =  REG_KEY_ID_W'('h205),
    CSR_VSSCRATCH      =  REG_KEY_ID_W'('h240),
    CSR_VSEPC          =  REG_KEY_ID_W'('h241),
    CSR_VSCAUSE        =  REG_KEY_ID_W'('h242),
    CSR_VSTVAL         =  REG_KEY_ID_W'('h243),
    CSR_VSIP           =  REG_KEY_ID_W'('h244),
    CSR_VSTIMECMP      =  REG_KEY_ID_W'('h24d),
    CSR_VSISELECT      =  REG_KEY_ID_W'('h250),
    CSR_VSIREG         =  REG_KEY_ID_W'('h251),
    CSR_VSIREG2        =  REG_KEY_ID_W'('h252),
    CSR_VSIREG3        =  REG_KEY_ID_W'('h253),
    CSR_VSIREG4        =  REG_KEY_ID_W'('h255),
    CSR_VSIREG5        =  REG_KEY_ID_W'('h256),
    CSR_VSIREG6        =  REG_KEY_ID_W'('h257),
    CSR_VSTOPEI        =  REG_KEY_ID_W'('h25c),
    CSR_VSATP          =  REG_KEY_ID_W'('h280),
    CSR_HSTATUS        =  REG_KEY_ID_W'('h600),
    CSR_HEDELEG        =  REG_KEY_ID_W'('h602),
    CSR_HIDELEG        =  REG_KEY_ID_W'('h603),
    CSR_HIE            =  REG_KEY_ID_W'('h604),
    CSR_HTIMEDELTA     =  REG_KEY_ID_W'('h605),
    CSR_HCOUNTEREN     =  REG_KEY_ID_W'('h606),
    CSR_HGEIE          =  REG_KEY_ID_W'('h607),
    CSR_HVIEN          =  REG_KEY_ID_W'('h608),
    CSR_HVICTL         =  REG_KEY_ID_W'('h609),
    CSR_HENVCFG        =  REG_KEY_ID_W'('h60a),
    CSR_HSTATEEN0      =  REG_KEY_ID_W'('h60c),
    CSR_HSTATEEN1      =  REG_KEY_ID_W'('h60d),
    CSR_HSTATEEN2      =  REG_KEY_ID_W'('h60e),
    CSR_HSTATEEN3      =  REG_KEY_ID_W'('h60f),
    CSR_HTVAL          =  REG_KEY_ID_W'('h643),
    CSR_HIP            =  REG_KEY_ID_W'('h644),
    CSR_HVIP           =  REG_KEY_ID_W'('h645),
    CSR_HVIPRIO1       =  REG_KEY_ID_W'('h646),
    CSR_HVIPRIO2       =  REG_KEY_ID_W'('h647),
    CSR_HTINST         =  REG_KEY_ID_W'('h64a),
    CSR_HGATP          =  REG_KEY_ID_W'('h680),
    CSR_HCONTEXT       =  REG_KEY_ID_W'('h6a8),
    CSR_HGEIP          =  REG_KEY_ID_W'('he12),
    CSR_VSTOPI         =  REG_KEY_ID_W'('heb0),
    CSR_SCOUNTOVF      =  REG_KEY_ID_W'('hda0),
    CSR_STOPI          =  REG_KEY_ID_W'('hdb0),
    CSR_UTVT           =  REG_KEY_ID_W'('h7),
    CSR_UNXTI          =  REG_KEY_ID_W'('h45),
    CSR_UINTSTATUS     =  REG_KEY_ID_W'('h46),
    CSR_USCRATCHCSW    =  REG_KEY_ID_W'('h48),
    CSR_USCRATCHCSWL   =  REG_KEY_ID_W'('h49),
    CSR_STVT           =  REG_KEY_ID_W'('h107),
    CSR_SNXTI          =  REG_KEY_ID_W'('h145),
    CSR_SINTSTATUS     =  REG_KEY_ID_W'('h146),
    CSR_SSCRATCHCSW    =  REG_KEY_ID_W'('h148),
    CSR_SSCRATCHCSWL   =  REG_KEY_ID_W'('h149),
    CSR_MTVT           =  REG_KEY_ID_W'('h307),
    CSR_MNXTI          =  REG_KEY_ID_W'('h345),
    CSR_MINTSTATUS     =  REG_KEY_ID_W'('h346),
    CSR_MSCRATCHCSW    =  REG_KEY_ID_W'('h348),
    CSR_MSCRATCHCSWL   =  REG_KEY_ID_W'('h349),
    CSR_MSTATUS        =  REG_KEY_ID_W'('h300),
    CSR_MISA           =  REG_KEY_ID_W'('h301),
    CSR_MEDELEG        =  REG_KEY_ID_W'('h302),
    CSR_MIDELEG        =  REG_KEY_ID_W'('h303),
    CSR_MIE            =  REG_KEY_ID_W'('h304),
    CSR_MTVEC          =  REG_KEY_ID_W'('h305),
    CSR_MCOUNTEREN     =  REG_KEY_ID_W'('h306),
    CSR_MVIEN          =  REG_KEY_ID_W'('h308),
    CSR_MVIP           =  REG_KEY_ID_W'('h309),
    CSR_MENVCFG        =  REG_KEY_ID_W'('h30a),
    CSR_MSTATEEN0      =  REG_KEY_ID_W'('h30c),
    CSR_MSTATEEN1      =  REG_KEY_ID_W'('h30d),
    CSR_MSTATEEN2      =  REG_KEY_ID_W'('h30e),
    CSR_MSTATEEN3      =  REG_KEY_ID_W'('h30f),
    CSR_MCOUNTINHIBIT  =  REG_KEY_ID_W'('h320),
    CSR_MSCRATCH       =  REG_KEY_ID_W'('h340),
    CSR_MEPC           =  REG_KEY_ID_W'('h341),
    CSR_MCAUSE         =  REG_KEY_ID_W'('h342),
    CSR_MTVAL          =  REG_KEY_ID_W'('h343),
    CSR_MIP            =  REG_KEY_ID_W'('h344),
    CSR_MTINST         =  REG_KEY_ID_W'('h34a),
    CSR_MTVAL2         =  REG_KEY_ID_W'('h34b),
    CSR_MISELECT       =  REG_KEY_ID_W'('h350),
    CSR_MIREG          =  REG_KEY_ID_W'('h351),
    CSR_MIREG2         =  REG_KEY_ID_W'('h352),
    CSR_MIREG3         =  REG_KEY_ID_W'('h353),
    CSR_MIREG4         =  REG_KEY_ID_W'('h355),
    CSR_MIREG5         =  REG_KEY_ID_W'('h356),
    CSR_MIREG6         =  REG_KEY_ID_W'('h357),
    CSR_MTOPEI         =  REG_KEY_ID_W'('h35c),
    CSR_PMPCFG0        =  REG_KEY_ID_W'('h3a0),
    CSR_PMPCFG1        =  REG_KEY_ID_W'('h3a1),
    CSR_PMPCFG2        =  REG_KEY_ID_W'('h3a2),
    CSR_PMPCFG3        =  REG_KEY_ID_W'('h3a3),
    CSR_PMPCFG4        =  REG_KEY_ID_W'('h3a4),
    CSR_PMPCFG5        =  REG_KEY_ID_W'('h3a5),
    CSR_PMPCFG6        =  REG_KEY_ID_W'('h3a6),
    CSR_PMPCFG7        =  REG_KEY_ID_W'('h3a7),
    CSR_PMPCFG8        =  REG_KEY_ID_W'('h3a8),
    CSR_PMPCFG9        =  REG_KEY_ID_W'('h3a9),
    CSR_PMPCFG10       =  REG_KEY_ID_W'('h3aa),
    CSR_PMPCFG11       =  REG_KEY_ID_W'('h3ab),
    CSR_PMPCFG12       =  REG_KEY_ID_W'('h3ac),
    CSR_PMPCFG13       =  REG_KEY_ID_W'('h3ad),
    CSR_PMPCFG14       =  REG_KEY_ID_W'('h3ae),
    CSR_PMPCFG15       =  REG_KEY_ID_W'('h3af),
    CSR_PMPADDR0       =  REG_KEY_ID_W'('h3b0),
    CSR_PMPADDR1       =  REG_KEY_ID_W'('h3b1),
    CSR_PMPADDR2       =  REG_KEY_ID_W'('h3b2),
    CSR_PMPADDR3       =  REG_KEY_ID_W'('h3b3),
    CSR_PMPADDR4       =  REG_KEY_ID_W'('h3b4),
    CSR_PMPADDR5       =  REG_KEY_ID_W'('h3b5),
    CSR_PMPADDR6       =  REG_KEY_ID_W'('h3b6),
    CSR_PMPADDR7       =  REG_KEY_ID_W'('h3b7),
    CSR_PMPADDR8       =  REG_KEY_ID_W'('h3b8),
    CSR_PMPADDR9       =  REG_KEY_ID_W'('h3b9),
    CSR_PMPADDR10      =  REG_KEY_ID_W'('h3ba),
    CSR_PMPADDR11      =  REG_KEY_ID_W'('h3bb),
    CSR_PMPADDR12      =  REG_KEY_ID_W'('h3bc),
    CSR_PMPADDR13      =  REG_KEY_ID_W'('h3bd),
    CSR_PMPADDR14      =  REG_KEY_ID_W'('h3be),
    CSR_PMPADDR15      =  REG_KEY_ID_W'('h3bf),
    CSR_PMPADDR16      =  REG_KEY_ID_W'('h3c0),
    CSR_PMPADDR17      =  REG_KEY_ID_W'('h3c1),
    CSR_PMPADDR18      =  REG_KEY_ID_W'('h3c2),
    CSR_PMPADDR19      =  REG_KEY_ID_W'('h3c3),
    CSR_PMPADDR20      =  REG_KEY_ID_W'('h3c4),
    CSR_PMPADDR21      =  REG_KEY_ID_W'('h3c5),
    CSR_PMPADDR22      =  REG_KEY_ID_W'('h3c6),
    CSR_PMPADDR23      =  REG_KEY_ID_W'('h3c7),
    CSR_PMPADDR24      =  REG_KEY_ID_W'('h3c8),
    CSR_PMPADDR25      =  REG_KEY_ID_W'('h3c9),
    CSR_PMPADDR26      =  REG_KEY_ID_W'('h3ca),
    CSR_PMPADDR27      =  REG_KEY_ID_W'('h3cb),
    CSR_PMPADDR28      =  REG_KEY_ID_W'('h3cc),
    CSR_PMPADDR29      =  REG_KEY_ID_W'('h3cd),
    CSR_PMPADDR30      =  REG_KEY_ID_W'('h3ce),
    CSR_PMPADDR31      =  REG_KEY_ID_W'('h3cf),
    CSR_PMPADDR32      =  REG_KEY_ID_W'('h3d0),
    CSR_PMPADDR33      =  REG_KEY_ID_W'('h3d1),
    CSR_PMPADDR34      =  REG_KEY_ID_W'('h3d2),
    CSR_PMPADDR35      =  REG_KEY_ID_W'('h3d3),
    CSR_PMPADDR36      =  REG_KEY_ID_W'('h3d4),
    CSR_PMPADDR37      =  REG_KEY_ID_W'('h3d5),
    CSR_PMPADDR38      =  REG_KEY_ID_W'('h3d6),
    CSR_PMPADDR39      =  REG_KEY_ID_W'('h3d7),
    CSR_PMPADDR40      =  REG_KEY_ID_W'('h3d8),
    CSR_PMPADDR41      =  REG_KEY_ID_W'('h3d9),
    CSR_PMPADDR42      =  REG_KEY_ID_W'('h3da),
    CSR_PMPADDR43      =  REG_KEY_ID_W'('h3db),
    CSR_PMPADDR44      =  REG_KEY_ID_W'('h3dc),
    CSR_PMPADDR45      =  REG_KEY_ID_W'('h3dd),
    CSR_PMPADDR46      =  REG_KEY_ID_W'('h3de),
    CSR_PMPADDR47      =  REG_KEY_ID_W'('h3df),
    CSR_PMPADDR48      =  REG_KEY_ID_W'('h3e0),
    CSR_PMPADDR49      =  REG_KEY_ID_W'('h3e1),
    CSR_PMPADDR50      =  REG_KEY_ID_W'('h3e2),
    CSR_PMPADDR51      =  REG_KEY_ID_W'('h3e3),
    CSR_PMPADDR52      =  REG_KEY_ID_W'('h3e4),
    CSR_PMPADDR53      =  REG_KEY_ID_W'('h3e5),
    CSR_PMPADDR54      =  REG_KEY_ID_W'('h3e6),
    CSR_PMPADDR55      =  REG_KEY_ID_W'('h3e7),
    CSR_PMPADDR56      =  REG_KEY_ID_W'('h3e8),
    CSR_PMPADDR57      =  REG_KEY_ID_W'('h3e9),
    CSR_PMPADDR58      =  REG_KEY_ID_W'('h3ea),
    CSR_PMPADDR59      =  REG_KEY_ID_W'('h3eb),
    CSR_PMPADDR60      =  REG_KEY_ID_W'('h3ec),
    CSR_PMPADDR61      =  REG_KEY_ID_W'('h3ed),
    CSR_PMPADDR62      =  REG_KEY_ID_W'('h3ee),
    CSR_PMPADDR63      =  REG_KEY_ID_W'('h3ef),
    CSR_MSECCFG        =  REG_KEY_ID_W'('h747),
    CSR_TSELECT        =  REG_KEY_ID_W'('h7a0),
    CSR_TDATA1         =  REG_KEY_ID_W'('h7a1),
    CSR_TDATA2         =  REG_KEY_ID_W'('h7a2),
    CSR_TDATA3         =  REG_KEY_ID_W'('h7a3),
    CSR_TINFO          =  REG_KEY_ID_W'('h7a4),
    CSR_TCONTROL       =  REG_KEY_ID_W'('h7a5),
    CSR_MCONTEXT       =  REG_KEY_ID_W'('h7a8),
    CSR_MSCONTEXT      =  REG_KEY_ID_W'('h7aa),
    CSR_DCSR           =  REG_KEY_ID_W'('h7b0),
    CSR_DPC            =  REG_KEY_ID_W'('h7b1),
    CSR_DSCRATCH0      =  REG_KEY_ID_W'('h7b2),
    CSR_DSCRATCH1      =  REG_KEY_ID_W'('h7b3),
    CSR_MCYCLE         =  REG_KEY_ID_W'('hb00),
    CSR_MINSTRET       =  REG_KEY_ID_W'('hb02),
    CSR_MHPMCOUNTER3   =  REG_KEY_ID_W'('hb03),
    CSR_MHPMCOUNTER4   =  REG_KEY_ID_W'('hb04),
    CSR_MHPMCOUNTER5   =  REG_KEY_ID_W'('hb05),
    CSR_MHPMCOUNTER6   =  REG_KEY_ID_W'('hb06),
    CSR_MHPMCOUNTER7   =  REG_KEY_ID_W'('hb07),
    CSR_MHPMCOUNTER8   =  REG_KEY_ID_W'('hb08),
    CSR_MHPMCOUNTER9   =  REG_KEY_ID_W'('hb09),
    CSR_MHPMCOUNTER10  =  REG_KEY_ID_W'('hb0a),
    CSR_MHPMCOUNTER11  =  REG_KEY_ID_W'('hb0b),
    CSR_MHPMCOUNTER12  =  REG_KEY_ID_W'('hb0c),
    CSR_MHPMCOUNTER13  =  REG_KEY_ID_W'('hb0d),
    CSR_MHPMCOUNTER14  =  REG_KEY_ID_W'('hb0e),
    CSR_MHPMCOUNTER15  =  REG_KEY_ID_W'('hb0f),
    CSR_MHPMCOUNTER16  =  REG_KEY_ID_W'('hb10),
    CSR_MHPMCOUNTER17  =  REG_KEY_ID_W'('hb11),
    CSR_MHPMCOUNTER18  =  REG_KEY_ID_W'('hb12),
    CSR_MHPMCOUNTER19  =  REG_KEY_ID_W'('hb13),
    CSR_MHPMCOUNTER20  =  REG_KEY_ID_W'('hb14),
    CSR_MHPMCOUNTER21  =  REG_KEY_ID_W'('hb15),
    CSR_MHPMCOUNTER22  =  REG_KEY_ID_W'('hb16),
    CSR_MHPMCOUNTER23  =  REG_KEY_ID_W'('hb17),
    CSR_MHPMCOUNTER24  =  REG_KEY_ID_W'('hb18),
    CSR_MHPMCOUNTER25  =  REG_KEY_ID_W'('hb19),
    CSR_MHPMCOUNTER26  =  REG_KEY_ID_W'('hb1a),
    CSR_MHPMCOUNTER27  =  REG_KEY_ID_W'('hb1b),
    CSR_MHPMCOUNTER28  =  REG_KEY_ID_W'('hb1c),
    CSR_MHPMCOUNTER29  =  REG_KEY_ID_W'('hb1d),
    CSR_MHPMCOUNTER30  =  REG_KEY_ID_W'('hb1e),
    CSR_MHPMCOUNTER31  =  REG_KEY_ID_W'('hb1f),
    CSR_MCYCLECFG      =  REG_KEY_ID_W'('h321),
    CSR_MINSTRETCFG    =  REG_KEY_ID_W'('h322),
    CSR_MHPMEVENT3     =  REG_KEY_ID_W'('h323),
    CSR_MHPMEVENT4     =  REG_KEY_ID_W'('h324),
    CSR_MHPMEVENT5     =  REG_KEY_ID_W'('h325),
    CSR_MHPMEVENT6     =  REG_KEY_ID_W'('h326),
    CSR_MHPMEVENT7     =  REG_KEY_ID_W'('h327),
    CSR_MHPMEVENT8     =  REG_KEY_ID_W'('h328),
    CSR_MHPMEVENT9     =  REG_KEY_ID_W'('h329),
    CSR_MHPMEVENT10    =  REG_KEY_ID_W'('h32a),
    CSR_MHPMEVENT11    =  REG_KEY_ID_W'('h32b),
    CSR_MHPMEVENT12    =  REG_KEY_ID_W'('h32c),
    CSR_MHPMEVENT13    =  REG_KEY_ID_W'('h32d),
    CSR_MHPMEVENT14    =  REG_KEY_ID_W'('h32e),
    CSR_MHPMEVENT15    =  REG_KEY_ID_W'('h32f),
    CSR_MHPMEVENT16    =  REG_KEY_ID_W'('h330),
    CSR_MHPMEVENT17    =  REG_KEY_ID_W'('h331),
    CSR_MHPMEVENT18    =  REG_KEY_ID_W'('h332),
    CSR_MHPMEVENT19    =  REG_KEY_ID_W'('h333),
    CSR_MHPMEVENT20    =  REG_KEY_ID_W'('h334),
    CSR_MHPMEVENT21    =  REG_KEY_ID_W'('h335),
    CSR_MHPMEVENT22    =  REG_KEY_ID_W'('h336),
    CSR_MHPMEVENT23    =  REG_KEY_ID_W'('h337),
    CSR_MHPMEVENT24    =  REG_KEY_ID_W'('h338),
    CSR_MHPMEVENT25    =  REG_KEY_ID_W'('h339),
    CSR_MHPMEVENT26    =  REG_KEY_ID_W'('h33a),
    CSR_MHPMEVENT27    =  REG_KEY_ID_W'('h33b),
    CSR_MHPMEVENT28    =  REG_KEY_ID_W'('h33c),
    CSR_MHPMEVENT29    =  REG_KEY_ID_W'('h33d),
    CSR_MHPMEVENT30    =  REG_KEY_ID_W'('h33e),
    CSR_MHPMEVENT31    =  REG_KEY_ID_W'('h33f),
    CSR_MVENDORID      =  REG_KEY_ID_W'('hf11),
    CSR_MARCHID        =  REG_KEY_ID_W'('hf12),
    CSR_MIMPID         =  REG_KEY_ID_W'('hf13),
    CSR_MHARTID        =  REG_KEY_ID_W'('hf14),
    CSR_MCONFIGPTR     =  REG_KEY_ID_W'('hf15),
    CSR_MTOPI          =  REG_KEY_ID_W'('hfb0),
    CSR_SIEH           =  REG_KEY_ID_W'('h114),
    CSR_SIPH           =  REG_KEY_ID_W'('h154),
    CSR_STIMECMPH      =  REG_KEY_ID_W'('h15d),
    CSR_VSIEH          =  REG_KEY_ID_W'('h214),
    CSR_VSIPH          =  REG_KEY_ID_W'('h254),
    CSR_VSTIMECMPH     =  REG_KEY_ID_W'('h25d),
    CSR_HTIMEDELTAH    =  REG_KEY_ID_W'('h615),
    CSR_HIDELEGH       =  REG_KEY_ID_W'('h613),
    CSR_HVIENH         =  REG_KEY_ID_W'('h618),
    CSR_HENVCFGH       =  REG_KEY_ID_W'('h61a),
    CSR_HVIPH          =  REG_KEY_ID_W'('h655),
    CSR_HVIPRIO1H      =  REG_KEY_ID_W'('h656),
    CSR_HVIPRIO2H      =  REG_KEY_ID_W'('h657),
    CSR_HSTATEEN0H     =  REG_KEY_ID_W'('h61c),
    CSR_HSTATEEN1H     =  REG_KEY_ID_W'('h61d),
    CSR_HSTATEEN2H     =  REG_KEY_ID_W'('h61e),
    CSR_HSTATEEN3H     =  REG_KEY_ID_W'('h61f),
    CSR_CYCLEH         =  REG_KEY_ID_W'('hc80),
    CSR_TIMEH          =  REG_KEY_ID_W'('hc81),
    CSR_INSTRETH       =  REG_KEY_ID_W'('hc82),
    CSR_HPMCOUNTER3H   =  REG_KEY_ID_W'('hc83),
    CSR_HPMCOUNTER4H   =  REG_KEY_ID_W'('hc84),
    CSR_HPMCOUNTER5H   =  REG_KEY_ID_W'('hc85),
    CSR_HPMCOUNTER6H   =  REG_KEY_ID_W'('hc86),
    CSR_HPMCOUNTER7H   =  REG_KEY_ID_W'('hc87),
    CSR_HPMCOUNTER8H   =  REG_KEY_ID_W'('hc88),
    CSR_HPMCOUNTER9H   =  REG_KEY_ID_W'('hc89),
    CSR_HPMCOUNTER10H  =  REG_KEY_ID_W'('hc8a),
    CSR_HPMCOUNTER11H  =  REG_KEY_ID_W'('hc8b),
    CSR_HPMCOUNTER12H  =  REG_KEY_ID_W'('hc8c),
    CSR_HPMCOUNTER13H  =  REG_KEY_ID_W'('hc8d),
    CSR_HPMCOUNTER14H  =  REG_KEY_ID_W'('hc8e),
    CSR_HPMCOUNTER15H  =  REG_KEY_ID_W'('hc8f),
    CSR_HPMCOUNTER16H  =  REG_KEY_ID_W'('hc90),
    CSR_HPMCOUNTER17H  =  REG_KEY_ID_W'('hc91),
    CSR_HPMCOUNTER18H  =  REG_KEY_ID_W'('hc92),
    CSR_HPMCOUNTER19H  =  REG_KEY_ID_W'('hc93),
    CSR_HPMCOUNTER20H  =  REG_KEY_ID_W'('hc94),
    CSR_HPMCOUNTER21H  =  REG_KEY_ID_W'('hc95),
    CSR_HPMCOUNTER22H  =  REG_KEY_ID_W'('hc96),
    CSR_HPMCOUNTER23H  =  REG_KEY_ID_W'('hc97),
    CSR_HPMCOUNTER24H  =  REG_KEY_ID_W'('hc98),
    CSR_HPMCOUNTER25H  =  REG_KEY_ID_W'('hc99),
    CSR_HPMCOUNTER26H  =  REG_KEY_ID_W'('hc9a),
    CSR_HPMCOUNTER27H  =  REG_KEY_ID_W'('hc9b),
    CSR_HPMCOUNTER28H  =  REG_KEY_ID_W'('hc9c),
    CSR_HPMCOUNTER29H  =  REG_KEY_ID_W'('hc9d),
    CSR_HPMCOUNTER30H  =  REG_KEY_ID_W'('hc9e),
    CSR_HPMCOUNTER31H  =  REG_KEY_ID_W'('hc9f),
    CSR_MSTATUSH       =  REG_KEY_ID_W'('h310),
    CSR_MIDELEGH       =  REG_KEY_ID_W'('h313),
    CSR_MIEH           =  REG_KEY_ID_W'('h314),
    CSR_MVIENH         =  REG_KEY_ID_W'('h318),
    CSR_MVIPH          =  REG_KEY_ID_W'('h319),
    CSR_MENVCFGH       =  REG_KEY_ID_W'('h31a),
    CSR_MSTATEEN0H     =  REG_KEY_ID_W'('h31c),
    CSR_MSTATEEN1H     =  REG_KEY_ID_W'('h31d),
    CSR_MSTATEEN2H     =  REG_KEY_ID_W'('h31e),
    CSR_MSTATEEN3H     =  REG_KEY_ID_W'('h31f),
    CSR_MIPH           =  REG_KEY_ID_W'('h354),
    CSR_MCYCLECFGH     =  REG_KEY_ID_W'('h721),
    CSR_MINSTRETCFGH   =  REG_KEY_ID_W'('h722),
    CSR_MHPMEVENT3H    =  REG_KEY_ID_W'('h723),
    CSR_MHPMEVENT4H    =  REG_KEY_ID_W'('h724),
    CSR_MHPMEVENT5H    =  REG_KEY_ID_W'('h725),
    CSR_MHPMEVENT6H    =  REG_KEY_ID_W'('h726),
    CSR_MHPMEVENT7H    =  REG_KEY_ID_W'('h727),
    CSR_MHPMEVENT8H    =  REG_KEY_ID_W'('h728),
    CSR_MHPMEVENT9H    =  REG_KEY_ID_W'('h729),
    CSR_MHPMEVENT10H   =  REG_KEY_ID_W'('h72a),
    CSR_MHPMEVENT11H   =  REG_KEY_ID_W'('h72b),
    CSR_MHPMEVENT12H   =  REG_KEY_ID_W'('h72c),
    CSR_MHPMEVENT13H   =  REG_KEY_ID_W'('h72d),
    CSR_MHPMEVENT14H   =  REG_KEY_ID_W'('h72e),
    CSR_MHPMEVENT15H   =  REG_KEY_ID_W'('h72f),
    CSR_MHPMEVENT16H   =  REG_KEY_ID_W'('h730),
    CSR_MHPMEVENT17H   =  REG_KEY_ID_W'('h731),
    CSR_MHPMEVENT18H   =  REG_KEY_ID_W'('h732),
    CSR_MHPMEVENT19H   =  REG_KEY_ID_W'('h733),
    CSR_MHPMEVENT20H   =  REG_KEY_ID_W'('h734),
    CSR_MHPMEVENT21H   =  REG_KEY_ID_W'('h735),
    CSR_MHPMEVENT22H   =  REG_KEY_ID_W'('h736),
    CSR_MHPMEVENT23H   =  REG_KEY_ID_W'('h737),
    CSR_MHPMEVENT24H   =  REG_KEY_ID_W'('h738),
    CSR_MHPMEVENT25H   =  REG_KEY_ID_W'('h739),
    CSR_MHPMEVENT26H   =  REG_KEY_ID_W'('h73a),
    CSR_MHPMEVENT27H   =  REG_KEY_ID_W'('h73b),
    CSR_MHPMEVENT28H   =  REG_KEY_ID_W'('h73c),
    CSR_MHPMEVENT29H   =  REG_KEY_ID_W'('h73d),
    CSR_MHPMEVENT30H   =  REG_KEY_ID_W'('h73e),
    CSR_MHPMEVENT31H   =  REG_KEY_ID_W'('h73f),
    CSR_MNSCRATCH      =  REG_KEY_ID_W'('h740),
    CSR_MNEPC          =  REG_KEY_ID_W'('h741),
    CSR_MNCAUSE        =  REG_KEY_ID_W'('h742),
    CSR_MNSTATUS       =  REG_KEY_ID_W'('h744),
    CSR_MSECCFGH       =  REG_KEY_ID_W'('h757),
    CSR_MCYCLEH        =  REG_KEY_ID_W'('hb80),
    CSR_MINSTRETH      =  REG_KEY_ID_W'('hb82),
    CSR_MHPMCOUNTER3H  =  REG_KEY_ID_W'('hb83),
    CSR_MHPMCOUNTER4H  =  REG_KEY_ID_W'('hb84),
    CSR_MHPMCOUNTER5H  =  REG_KEY_ID_W'('hb85),
    CSR_MHPMCOUNTER6H  =  REG_KEY_ID_W'('hb86),
    CSR_MHPMCOUNTER7H  =  REG_KEY_ID_W'('hb87),
    CSR_MHPMCOUNTER8H  =  REG_KEY_ID_W'('hb88),
    CSR_MHPMCOUNTER9H  =  REG_KEY_ID_W'('hb89),
    CSR_MHPMCOUNTER10H =  REG_KEY_ID_W'('hb8a),
    CSR_MHPMCOUNTER11H =  REG_KEY_ID_W'('hb8b),
    CSR_MHPMCOUNTER12H =  REG_KEY_ID_W'('hb8c),
    CSR_MHPMCOUNTER13H =  REG_KEY_ID_W'('hb8d),
    CSR_MHPMCOUNTER14H =  REG_KEY_ID_W'('hb8e),
    CSR_MHPMCOUNTER15H =  REG_KEY_ID_W'('hb8f),
    CSR_MHPMCOUNTER16H =  REG_KEY_ID_W'('hb90),
    CSR_MHPMCOUNTER17H =  REG_KEY_ID_W'('hb91),
    CSR_MHPMCOUNTER18H =  REG_KEY_ID_W'('hb92),
    CSR_MHPMCOUNTER19H =  REG_KEY_ID_W'('hb93),
    CSR_MHPMCOUNTER20H =  REG_KEY_ID_W'('hb94),
    CSR_MHPMCOUNTER21H =  REG_KEY_ID_W'('hb95),
    CSR_MHPMCOUNTER22H =  REG_KEY_ID_W'('hb96),
    CSR_MHPMCOUNTER23H =  REG_KEY_ID_W'('hb97),
    CSR_MHPMCOUNTER24H =  REG_KEY_ID_W'('hb98),
    CSR_MHPMCOUNTER25H =  REG_KEY_ID_W'('hb99),
    CSR_MHPMCOUNTER26H =  REG_KEY_ID_W'('hb9a),
    CSR_MHPMCOUNTER27H =  REG_KEY_ID_W'('hb9b),
    CSR_MHPMCOUNTER28H =  REG_KEY_ID_W'('hb9c),
    CSR_MHPMCOUNTER29H =  REG_KEY_ID_W'('hb9d),
    CSR_MHPMCOUNTER30H =  REG_KEY_ID_W'('hb9e),
    CSR_MHPMCOUNTER31H =  REG_KEY_ID_W'('hb9f)
  } csr_id_e;
endpackage